library verilog;
use verilog.vl_types.all;
entity clockDivider_testbench is
end clockDivider_testbench;
